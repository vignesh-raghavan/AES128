module isbox (
	input [7:0] index,

	output [7:0] o
);

wire a, b, c, d, e, f, g, h;

assign a = index[7];
assign b = index[6];
assign c = index[5];
assign d = index[4];
assign e = index[3];
assign f = index[2];
assign g = index[1];
assign h = index[0];


wire [620:0] x;



assign x[0] = ( a & b & (~c) & d & (~e) & (~f) & g & h );
assign x[1] = ( a & (~c) & (~d) & e & f & (~g) & h );
assign x[2] = ( (~a) & (~b) & c & d & (~e) & (~f) & g & (~h) );
assign x[3] = ( (~a) & (~b) & c & d & (~e) & f & g & h );
assign x[4] = ( (~a) & (~b) & c & d & e & (~f) & g & (~h) );
assign x[5] = ( a & b & (~c) & (~d) & (~e) & (~f) & g & (~h) );
assign x[6] = ( (~a) & b & (~c) & d & (~e) & f & g & h );
assign x[7] = ( a & b & (~c) & d & e & (~f) & g & h );
assign x[8] = ( (~a) & b & c & d & e & f & g & (~h) );
assign x[9] = ( (~a) & (~b) & c & (~d) & (~e) & f & (~g) & (~h) );
assign x[10] = ( a & b & c & d & (~e) & f & (~g) & (~h) );
assign x[11] = ( a & b & (~c) & d & (~e) & f & (~g) & h );
assign x[12] = ( (~a) & b & (~c) & (~d) & (~e) & f & (~g) & (~h) );
assign x[13] = ( a & b & (~c) & d & e & (~f) & (~g) & h );
assign x[14] = ( (~a) & (~c) & (~d) & e & (~f) & g & h );
assign x[15] = ( (~a) & b & c & (~d) & (~f) & (~g) & (~h) );
assign x[16] = ( (~a) & b & (~c) & (~d) & (~e) & g & (~h) );
assign x[17] = ( a & (~b) & c & d & e & (~f) & g );
assign x[18] = ( (~a) & b & (~c) & (~e) & f & g & (~h) );
assign x[19] = ( (~a) & (~b) & (~c) & d & (~e) & g & h );
assign x[20] = ( (~a) & b & c & d & (~e) & (~g) & (~h) );
assign x[21] = ( a & (~b) & (~d) & (~e) & f & g & h );
assign x[22] = ( a & (~b) & c & d & e & (~f) & (~g) );
assign x[23] = ( a & b & c & (~d) & (~e) & (~g) & (~h) );
assign x[24] = ( a & (~c) & d & e & f & g & (~h) );
assign x[25] = ( a & b & (~d) & (~e) & f & (~g) & (~h) );
assign x[26] = ( a & c & (~d) & e & f & (~g) & (~h) );
assign x[27] = ( (~a) & (~b) & c & d & e & f & g & (~h) );
assign x[28] = ( a & b & c & d & e & (~f) & (~g) & (~h) );
assign x[29] = ( a & (~b) & (~c) & d & (~e) & (~f) & (~g) & (~h) );
assign x[30] = ( a & (~b) & (~c) & (~d) & e & f & (~g) & (~h) );
assign x[31] = ( a & (~b) & (~c) & d & e & (~f) & (~g) & (~h) );
assign x[32] = ( a & b & (~c) & d & e & f & (~g) & (~h) );
assign x[33] = ( b & (~d) & e & (~f) & (~g) & (~h) );
assign x[34] = ( (~a) & (~b) & c & (~d) & (~f) & g & (~h) );
assign x[35] = ( (~a) & (~b) & (~c) & (~d) & (~f) & g & h );
assign x[36] = ( (~a) & b & c & e & (~f) & (~g) & (~h) );
assign x[37] = ( a & b & c & (~d) & e & g & (~h) );
assign x[38] = ( a & b & c & (~d) & (~e) & f & g );
assign x[39] = ( a & b & c & (~e) & f & g & (~h) );
assign x[40] = ( (~a) & (~b) & c & (~d) & f & (~g) & h );
assign x[41] = ( (~a) & (~b) & (~c) & (~d) & f & g & (~h) );
assign x[42] = ( (~b) & c & d & (~e) & f & (~g) & h );
assign x[43] = ( (~a) & c & (~d) & e & (~f) & (~g) & (~h) );
assign x[44] = ( (~b) & (~c) & d & (~e) & f & g & h );
assign x[45] = ( b & c & (~d) & (~e) & f & (~g) & (~h) );
assign x[46] = ( (~a) & (~b) & (~c) & d & (~e) & f & (~h) );
assign x[47] = ( a & b & (~c) & d & e & f & h );
assign x[48] = ( (~a) & (~b) & (~c) & d & e & f & (~g) );
assign x[49] = ( (~a) & (~b) & d & e & f & (~g) & h );
assign x[50] = ( (~a) & b & c & (~d) & (~e) & (~f) & g & (~h) );
assign x[51] = ( (~a) & b & c & d & (~e) & (~f) & g & h );
assign x[52] = ( (~a) & b & c & (~d) & (~e) & f & (~g) & h );
assign x[53] = ( (~a) & (~b) & (~c) & d & (~e) & (~f) & (~g) & h );
assign x[54] = ( (~a) & b & c & d & e & (~f) & (~g) & h );
assign x[55] = ( a & (~b) & c & d & e & f & (~g) & h );
assign x[56] = ( (~a) & b & (~c) & d & e & f & (~g) & (~h) );
assign x[57] = ( (~a) & b & c & (~d) & e & (~g) );
assign x[58] = ( (~a) & (~b) & (~d) & e & g & (~h) );
assign x[59] = ( (~a) & (~b) & (~c) & (~d) & e & f );
assign x[60] = ( a & c & (~d) & (~f) & (~g) & h );
assign x[61] = ( b & (~d) & (~e) & (~f) & (~g) & h );
assign x[62] = ( a & (~b) & (~d) & (~f) & (~g) & h );
assign x[63] = ( (~a) & b & (~d) & e & (~f) & (~g) );
assign x[64] = ( b & (~c) & d & e & f & g );
assign x[65] = ( b & c & (~d) & (~e) & f & g & (~h) );
assign x[66] = ( a & (~b) & c & d & e & g & h );
assign x[67] = ( (~a) & (~b) & (~c) & d & f & g & (~h) );
assign x[68] = ( a & (~b) & (~c) & d & e & (~f) & h );
assign x[69] = ( (~a) & b & (~c) & d & f & (~g) & h );
assign x[70] = ( (~a) & (~b) & (~c) & d & e & (~g) & h );
assign x[71] = ( a & (~b) & (~c) & d & (~e) & (~g) & h );
assign x[72] = ( (~a) & b & (~c) & d & (~e) & f & (~g) );
assign x[73] = ( a & (~c) & (~d) & e & f & g & (~h) );
assign x[74] = ( (~a) & b & c & d & e & (~f) & g & (~h) );
assign x[75] = ( a & (~b) & d & (~e) & f & (~g) & (~h) );
assign x[76] = ( a & (~b) & c & d & (~e) & (~f) & (~g) & (~h) );
assign x[77] = ( a & (~b) & c & (~d) & e & f & g & (~h) );
assign x[78] = ( (~a) & (~c) & (~d) & e & f & g );
assign x[79] = ( a & (~d) & (~e) & f & g & (~h) );
assign x[80] = ( (~a) & (~b) & (~c) & e & f & g & h );
assign x[81] = ( a & (~b) & (~c) & (~d) & e & (~f) & g );
assign x[82] = ( (~b) & (~c) & (~d) & e & (~f) & (~g) & (~h) );


assign o[7] = |(x[82:0]);



assign x[83] = ( a & b & c & (~d) & e & (~g) & h );
assign x[84] = ( (~b) & (~c) & (~d) & e & (~f) & (~g) & h );
assign x[85] = ( (~a) & (~b) & c & (~d) & (~e) & (~f) & (~g) & (~h) );
assign x[86] = ( (~a) & b & c & (~d) & e & f & g & (~h) );
assign x[87] = ( (~a) & (~b) & (~c) & d & e & (~f) & g & (~h) );
assign x[88] = ( (~a) & c & (~d) & (~e) & (~f) & (~g) & h );
assign x[89] = ( (~b) & (~c) & (~d) & (~e) & (~f) & g & h );
assign x[90] = ( (~a) & (~b) & c & d & e & (~f) & h );
assign x[91] = ( (~a) & b & (~c) & d & (~e) & g & h );
assign x[92] = ( (~a) & (~c) & d & e & (~f) & g & h );
assign x[93] = ( b & (~c) & d & (~e) & (~f) & g & (~h) );
assign x[94] = ( x[17] );
assign x[95] = ( x[20] );
assign x[96] = ( b & (~c) & d & (~e) & (~f) & (~g) & (~h) );
assign x[97] = ( (~b) & (~c) & d & e & f & (~g) & h );
assign x[98] = ( a & c & d & e & f & (~g) & (~h) );
assign x[99] = ( a & b & c & (~d) & (~e) & (~f) & g & h );
assign x[100] = ( a & (~b) & c & d & (~e) & (~f) & g & h );
assign x[101] = ( a & b & c & d & (~e) & (~f) & g & h );
assign x[102] = ( (~a) & (~b) & c & d & (~e) & (~f) & g & h );
assign x[103] = ( a & (~b) & c & d & (~e) & (~f) & (~g) & h );
assign x[104] = ( x[27] );
assign x[105] = ( x[28] );
assign x[106] = ( x[30] );
assign x[107] = ( x[31] );
assign x[108] = ( b & c & (~d) & e & (~f) & (~g) );
assign x[109] = ( (~a) & b & (~c) & (~e) & (~f) & (~g) & h );
assign x[110] = ( (~a) & (~b) & c & (~d) & e & (~f) & (~g) );
assign x[111] = ( a & b & (~c) & (~e) & (~f) & (~g) & h );
assign x[112] = ( a & b & c & e & f & g & h );
assign x[113] = ( (~a) & b & (~c) & (~e) & f & (~g) & h );
assign x[114] = ( x[36] );
assign x[115] = ( a & c & d & e & (~f) & g & h );
assign x[116] = ( x[39] );
assign x[117] = ( a & (~b) & c & (~d) & e & (~f) & (~h) );
assign x[118] = ( (~a) & b & (~c) & (~d) & e & f & (~g) );
assign x[119] = ( a & (~c) & d & (~e) & (~f) & g & (~h) );
assign x[120] = ( x[40] );
assign x[121] = ( a & (~b) & (~c) & (~d) & f & g & h );
assign x[122] = ( (~a) & (~b) & c & d & e & (~g) & (~h) );
assign x[123] = ( a & c & d & (~e) & f & (~g) & h );
assign x[124] = ( x[42] );
assign x[125] = ( a & b & (~c) & d & (~e) & g & (~h) );
assign x[126] = ( (~a) & (~b) & (~d) & e & f & (~g) & h );
assign x[127] = ( (~a) & b & (~c) & d & e & (~f) & (~h) );
assign x[128] = ( x[47] );
assign x[129] = ( x[48] );
assign x[130] = ( (~a) & b & c & d & e & f & g & h );
assign x[131] = ( a & (~b) & c & d & (~e) & f & g & (~h) );
assign x[132] = ( x[53] );
assign x[133] = ( x[55] );
assign x[134] = ( (~a) & b & (~c) & (~d) & (~f) & g );
assign x[135] = ( (~a) & (~b) & c & (~d) & e & f );
assign x[136] = ( (~a) & b & (~d) & e & (~f) & (~h) );
assign x[137] = ( (~a) & (~c) & (~d) & (~e) & (~f) & (~h) );
assign x[138] = ( (~b) & (~c) & (~d) & e & f & g );
assign x[139] = ( x[61] );
assign x[140] = ( a & d & e & (~f) & (~g) & h );
assign x[141] = ( a & (~b) & c & (~d) & (~e) & (~f) & h );
assign x[142] = ( a & b & (~c) & (~d) & e & g & h );
assign x[143] = ( x[65] );
assign x[144] = ( a & (~b) & c & (~d) & (~f) & (~g) & (~h) );
assign x[145] = ( x[66] );
assign x[146] = ( (~a) & (~c) & d & (~e) & (~f) & (~g) & (~h) );
assign x[147] = ( a & (~b) & (~c) & (~d) & (~e) & f & (~g) );
assign x[148] = ( a & b & (~c) & d & (~f) & g & (~h) );
assign x[149] = ( x[67] );
assign x[150] = ( x[68] );
assign x[151] = ( a & (~b) & d & e & f & g & (~h) );
assign x[152] = ( x[72] );
assign x[153] = ( x[73] );
assign x[154] = ( x[75] );
assign x[155] = ( x[76] );
assign x[156] = ( x[79] );
assign x[157] = ( x[80] );
assign x[158] = ( x[81] );
assign x[159] = ( a & (~c) & d & e & f & g & h );


assign o[6] = |(x[159:83]);



assign x[160] = ( a & (~b) & (~c) & d & (~e) & (~f) & g & h );
assign x[161] = ( a & (~b) & (~c) & (~d) & (~e) & (~f) & (~g) & (~h) );
assign x[162] = ( a & b & (~c) & d & (~e) & (~f) & g & h );
assign x[163] = ( (~a) & (~c) & d & (~e) & f & g & (~h) );
assign x[164] = ( x[2] );
assign x[165] = ( a & b & (~c) & (~d) & e & (~f) & (~g) & (~h) );
assign x[166] = ( x[4] );
assign x[167] = ( x[5] );
assign x[168] = ( x[10] );
assign x[169] = ( x[11] );
assign x[170] = ( x[13] );
assign x[171] = ( (~a) & (~b) & (~c) & (~e) & (~f) & g & (~h) );
assign x[172] = ( (~a) & b & c & d & (~e) & (~g) & h );
assign x[173] = ( (~a) & (~b) & (~c) & (~d) & e & (~f) & (~h) );
assign x[174] = ( (~a) & (~b) & c & d & f & (~g) & (~h) );
assign x[175] = ( a & (~b) & (~d) & (~e) & f & (~g) & h );
assign x[176] = ( a & (~b) & c & e & f & (~g) & (~h) );
assign x[177] = ( a & (~b) & d & (~e) & (~f) & g & (~h) );
assign x[178] = ( (~a) & (~b) & d & (~e) & f & g & (~h) );
assign x[179] = ( x[23] );
assign x[180] = ( x[96] );
assign x[181] = ( b & (~c) & (~d) & e & f & g & (~h) );
assign x[182] = ( a & b & (~c) & (~d) & e & f & (~h) );
assign x[183] = ( a & b & c & (~d) & e & (~f) & g & h );
assign x[184] = ( x[102] );
assign x[185] = ( (~a) & (~b) & c & d & (~e) & (~f) & (~g) & h );
assign x[186] = ( x[28] );
assign x[187] = ( a & b & (~c) & d & e & (~f) & (~g) & (~h) );
assign x[188] = ( x[30] );
assign x[189] = ( x[31] );
assign x[190] = ( (~a) & b & (~c) & (~d) & (~e) & (~f) );
assign x[191] = ( (~b) & c & d & f & g & h );
assign x[192] = ( (~a) & b & (~d) & e & (~g) & h );
assign x[193] = ( (~a) & (~b) & (~d) & (~e) & f & (~h) );
assign x[194] = ( (~a) & (~b) & c & (~d) & (~e) & (~f) & h );
assign x[195] = ( x[109] );
assign x[196] = ( a & b & (~c) & (~d) & (~e) & g & h );
assign x[197] = ( (~a) & (~b) & (~d) & (~e) & f & g & h );
assign x[198] = ( x[112] );
assign x[199] = ( x[113] );
assign x[200] = ( x[38] );
assign x[201] = ( (~a) & (~b) & (~c) & e & (~f) & (~g) & (~h) );
assign x[202] = ( x[115] );
assign x[203] = ( x[117] );
assign x[204] = ( a & b & c & (~d) & (~e) & f & (~g) );
assign x[205] = ( (~a) & (~b) & (~c) & (~e) & f & (~g) & h );
assign x[206] = ( x[121] );
assign x[207] = ( x[122] );
assign x[208] = ( x[43] );
assign x[209] = ( x[126] );
assign x[210] = ( a & (~b) & (~c) & d & (~e) & f & (~h) );
assign x[211] = ( x[50] );
assign x[212] = ( x[130] );
assign x[213] = ( x[131] );
assign x[214] = ( x[52] );
assign x[215] = ( x[53] );
assign x[216] = ( x[54] );
assign x[217] = ( a & (~b) & (~c) & d & e & (~f) & g & (~h) );
assign x[218] = ( x[56] );
assign x[219] = ( (~a) & (~b) & (~c) & (~d) & f & h );
assign x[220] = ( a & b & c & d & (~g) & h );
assign x[221] = ( a & (~b) & (~c) & e & (~g) & h );
assign x[222] = ( a & b & c & d & (~e) & h );
assign x[223] = ( x[57] );
assign x[224] = ( x[60] );
assign x[225] = ( x[141] );
assign x[226] = ( x[146] );
assign x[227] = ( x[148] );
assign x[228] = ( x[67] );
assign x[229] = ( x[68] );
assign x[230] = ( x[71] );
assign x[231] = ( x[72] );
assign x[232] = ( x[73] );
assign x[233] = ( x[74] );
assign x[234] = ( x[76] );
assign x[235] = ( x[77] );
assign x[236] = ( a & b & c & (~d) & (~f) & g & (~h) );
assign x[237] = ( x[159] );


assign o[5] = |(x[237:160]);



assign x[238] = ( (~a) & b & (~c) & d & e & (~f) & (~g) & (~h) );
assign x[239] = ( (~a) & b & c & d & (~e) & (~f) & (~h) );
assign x[240] = ( x[85] );
assign x[241] = ( (~a) & b & (~c) & (~d) & (~e) & f & g & h );
assign x[242] = ( x[3] );
assign x[243] = ( a & b & c & d & e & f & g & h );
assign x[244] = ( x[165] );
assign x[245] = ( x[7] );
assign x[246] = ( x[10] );
assign x[247] = ( x[11] );
assign x[248] = ( x[88] );
assign x[249] = ( x[91] );
assign x[250] = ( (~a) & (~b) & (~c) & d & (~e) & g & (~h) );
assign x[251] = ( (~b) & c & (~d) & e & f & (~g) & h );
assign x[252] = ( x[15] );
assign x[253] = ( x[16] );
assign x[254] = ( (~a) & b & c & d & f & (~g) & h );
assign x[255] = ( a & (~c) & (~d) & e & (~f) & (~g) & h );
assign x[256] = ( (~a) & b & (~d) & e & f & (~g) & (~h) );
assign x[257] = ( b & (~c) & d & (~e) & f & (~g) & (~h) );
assign x[258] = ( x[97] );
assign x[259] = ( x[98] );
assign x[260] = ( x[101] );
assign x[261] = ( x[183] );
assign x[262] = ( x[24] );
assign x[263] = ( a & (~b) & c & (~d) & (~e) & f & (~g) & (~h) );
assign x[264] = ( x[103] );
assign x[265] = ( x[27] );
assign x[266] = ( a & b & c & d & (~e) & (~f) & (~g) & (~h) );
assign x[267] = ( x[29] );
assign x[268] = ( x[30] );
assign x[269] = ( x[32] );
assign x[270] = ( (~a) & (~b) & (~c) & (~e) & (~g) & (~h) );
assign x[271] = ( a & (~b) & (~c) & (~e) & g & (~h) );
assign x[272] = ( a & b & e & (~f) & g & (~h) );
assign x[273] = ( x[194] );
assign x[274] = ( a & (~b) & c & (~e) & (~f) & g & (~h) );
assign x[275] = ( x[109] );
assign x[276] = ( x[196] );
assign x[277] = ( x[197] );
assign x[278] = ( x[111] );
assign x[279] = ( x[34] );
assign x[280] = ( x[35] );
assign x[281] = ( (~a) & b & (~c) & d & e & (~f) & h );
assign x[282] = ( (~a) & b & (~c) & d & f & g & (~h) );
assign x[283] = ( b & c & (~d) & e & f & (~g) & h );
assign x[284] = ( x[37] );
assign x[285] = ( x[38] );
assign x[286] = ( x[201] );
assign x[287] = ( a & (~b) & (~d) & e & f & g & h );
assign x[288] = ( x[39] );
assign x[289] = ( x[119] );
assign x[290] = ( x[123] );
assign x[291] = ( x[42] );
assign x[292] = ( a & (~b) & (~c) & d & e & f & (~h) );
assign x[293] = ( x[131] );
assign x[294] = ( x[52] );
assign x[295] = ( x[217] );
assign x[296] = ( x[219] );
assign x[297] = ( x[136] );
assign x[298] = ( (~b) & c & d & e & (~f) & (~g) );
assign x[299] = ( x[221] );
assign x[300] = ( (~c) & (~d) & (~e) & (~f) & (~g) & (~h) );
assign x[301] = ( x[62] );
assign x[302] = ( x[141] );
assign x[303] = ( x[142] );
assign x[304] = ( x[65] );
assign x[305] = ( x[66] );
assign x[306] = ( x[151] );
assign x[307] = ( x[74] );
assign x[308] = ( x[76] );
assign x[309] = ( x[77] );
assign x[310] = ( x[78] );
assign x[311] = ( x[236] );
assign x[312] = ( x[82] );


assign o[4] = |(x[312:238]);



assign x[313] = ( (~a) & b & c & (~d) & (~e) & f & g & h );
assign x[314] = ( x[161] );
assign x[315] = ( x[238] );
assign x[316] = ( (~a) & b & (~d) & e & (~f) & g & (~h) );
assign x[317] = ( a & c & (~d) & e & (~f) & (~g) & (~h) );
assign x[318] = ( (~a) & (~b) & (~d) & e & (~f) & (~g) & (~h) );
assign x[319] = ( a & (~b) & (~c) & (~d) & (~e) & f & (~h) );
assign x[320] = ( a & b & c & (~d) & e & (~f) & (~g) & h );
assign x[321] = ( x[243] );
assign x[322] = ( x[5] );
assign x[323] = ( x[6] );
assign x[324] = ( x[8] );
assign x[325] = ( x[171] );
assign x[326] = ( (~a) & (~b) & c & (~d) & f & g & h );
assign x[327] = ( x[251] );
assign x[328] = ( x[14] );
assign x[329] = ( x[93] );
assign x[330] = ( x[18] );
assign x[331] = ( x[174] );
assign x[332] = ( x[176] );
assign x[333] = ( x[21] );
assign x[334] = ( x[256] );
assign x[335] = ( x[22] );
assign x[336] = ( x[99] );
assign x[337] = ( x[100] );
assign x[338] = ( x[101] );
assign x[339] = ( x[183] );
assign x[340] = ( x[25] );
assign x[341] = ( x[185] );
assign x[342] = ( x[263] );
assign x[343] = ( x[187] );
assign x[344] = ( (~a) & (~d) & (~e) & (~f) & (~g) & h );
assign x[345] = ( (~b) & c & d & e & (~f) & h );
assign x[346] = ( a & (~b) & c & (~d) & f & h );
assign x[347] = ( b & c & d & (~f) & (~g) & h );
assign x[348] = ( (~a) & (~b) & d & (~e) & (~g) & (~h) );
assign x[349] = ( a & b & e & f & g & (~h) );
assign x[350] = ( b & d & (~e) & f & (~g) & (~h) );
assign x[351] = ( x[274] );
assign x[352] = ( x[197] );
assign x[353] = ( x[110] );
assign x[354] = ( (~a) & b & c & d & (~e) & g & (~h) );
assign x[355] = ( x[113] );
assign x[356] = ( x[282] );
assign x[357] = ( a & b & (~c) & (~d) & (~e) & (~f) & (~g) );
assign x[358] = ( x[204] );
assign x[359] = ( x[125] );
assign x[360] = ( x[45] );
assign x[361] = ( x[292] );
assign x[362] = ( x[47] );
assign x[363] = ( x[49] );
assign x[364] = ( x[50] );
assign x[365] = ( x[51] );
assign x[366] = ( x[130] );
assign x[367] = ( x[131] );
assign x[368] = ( x[52] );
assign x[369] = ( x[55] );
assign x[370] = ( (~b) & (~d) & e & (~f) & g & h );
assign x[371] = ( a & b & (~c) & d & g & h );
assign x[372] = ( (~a) & d & (~e) & f & (~g) & h );
assign x[373] = ( x[142] );
assign x[374] = ( x[146] );
assign x[375] = ( x[148] );
assign x[376] = ( x[67] );
assign x[377] = ( x[68] );
assign x[378] = ( x[69] );
assign x[379] = ( x[151] );
assign x[380] = ( x[70] );
assign x[381] = ( x[71] );
assign x[382] = ( x[74] );
assign x[383] = ( x[76] );
assign x[384] = ( x[77] );
assign x[385] = ( x[236] );
assign x[386] = ( x[80] );
assign x[387] = ( x[81] );
assign x[388] = ( x[159] );


assign o[3] = |(x[388:313]);



assign x[389] = ( (~a) & (~b) & c & d & e & f & g & h );
assign x[390] = ( a & b & c & d & e & f & (~g) & (~h) );
assign x[391] = ( a & (~b) & c & (~d) & e & (~f) & h );
assign x[392] = ( x[85] );
assign x[393] = ( x[86] );
assign x[394] = ( x[241] );
assign x[395] = ( x[243] );
assign x[396] = ( x[7] );
assign x[397] = ( x[9] );
assign x[398] = ( x[12] );
assign x[399] = ( x[13] );
assign x[400] = ( x[326] );
assign x[401] = ( (~a) & c & (~d) & e & f & g & h );
assign x[402] = ( x[172] );
assign x[403] = ( x[92] );
assign x[404] = ( a & b & (~c) & e & f & g & h );
assign x[405] = ( x[177] );
assign x[406] = ( x[178] );
assign x[407] = ( x[181] );
assign x[408] = ( x[99] );
assign x[409] = ( x[182] );
assign x[410] = ( x[101] );
assign x[411] = ( x[183] );
assign x[412] = ( x[102] );
assign x[413] = ( x[185] );
assign x[414] = ( x[263] );
assign x[415] = ( x[103] );
assign x[416] = ( x[266] );
assign x[417] = ( x[187] );
assign x[418] = ( x[29] );
assign x[419] = ( (~a) & b & (~d) & e & (~f) & h );
assign x[420] = ( a & b & c & d & g & (~h) );
assign x[421] = ( a & (~b) & (~c) & f & (~g) & h );
assign x[422] = ( a & b & d & (~e) & f & h );
assign x[423] = ( x[110] );
assign x[424] = ( x[34] );
assign x[425] = ( x[35] );
assign x[426] = ( x[281] );
assign x[427] = ( x[354] );
assign x[428] = ( x[357] );
assign x[429] = ( x[201] );
assign x[430] = ( x[205] );
assign x[431] = ( x[118] );
assign x[432] = ( x[119] );
assign x[433] = ( x[122] );
assign x[434] = ( x[41] );
assign x[435] = ( x[44] );
assign x[436] = ( a & (~c) & (~d) & (~e) & f & (~g) & h );
assign x[437] = ( x[127] );
assign x[438] = ( x[45] );
assign x[439] = ( x[210] );
assign x[440] = ( x[292] );
assign x[441] = ( x[48] );
assign x[442] = ( x[51] );
assign x[443] = ( x[52] );
assign x[444] = ( x[54] );
assign x[445] = ( x[217] );
assign x[446] = ( x[55] );
assign x[447] = ( x[56] );
assign x[448] = ( x[134] );
assign x[449] = ( x[63] );
assign x[450] = ( x[64] );
assign x[451] = ( x[144] );
assign x[452] = ( x[66] );
assign x[453] = ( x[146] );
assign x[454] = ( x[147] );
assign x[455] = ( x[69] );
assign x[456] = ( x[70] );
assign x[457] = ( x[71] );
assign x[458] = ( x[72] );
assign x[459] = ( x[73] );
assign x[460] = ( x[74] );
assign x[461] = ( x[75] );
assign x[462] = ( x[76] );
assign x[463] = ( x[77] );
assign x[464] = ( x[79] );
assign x[465] = ( x[81] );
assign x[466] = ( x[82] );
assign x[467] = ( x[159] );


assign o[2] = |(x[467:389]);



assign x[468] = ( a & b & (~c) & (~d) & (~e) & (~f) & g & h );
assign x[469] = ( x[313] );
assign x[470] = ( x[160] );
assign x[471] = ( a & b & (~c) & (~d) & (~e) & f & g & (~h) );
assign x[472] = ( (~a) & c & (~d) & (~e) & f & g & (~h) );
assign x[473] = ( x[320] );
assign x[474] = ( x[241] );
assign x[475] = ( x[3] );
assign x[476] = ( x[87] );
assign x[477] = ( x[4] );
assign x[478] = ( x[6] );
assign x[479] = ( x[8] );
assign x[480] = ( x[9] );
assign x[481] = ( x[12] );
assign x[482] = ( a & (~b) & c & e & (~f) & (~g) & h );
assign x[483] = ( x[401] );
assign x[484] = ( x[254] );
assign x[485] = ( x[173] );
assign x[486] = ( x[19] );
assign x[487] = ( x[255] );
assign x[488] = ( x[404] );
assign x[489] = ( a & b & (~d) & e & f & (~g) & (~h) );
assign x[490] = ( x[100] );
assign x[491] = ( x[102] );
assign x[492] = ( x[26] );
assign x[493] = ( x[185] );
assign x[494] = ( x[103] );
assign x[495] = ( x[266] );
assign x[496] = ( x[29] );
assign x[497] = ( x[31] );
assign x[498] = ( x[32] );
assign x[499] = ( x[194] );
assign x[500] = ( x[274] );
assign x[501] = ( x[354] );
assign x[502] = ( x[283] );
assign x[503] = ( x[115] );
assign x[504] = ( x[287] );
assign x[505] = ( x[117] );
assign x[506] = ( x[204] );
assign x[507] = ( x[205] );
assign x[508] = ( x[40] );
assign x[509] = ( x[121] );
assign x[510] = ( x[123] );
assign x[511] = ( x[125] );
assign x[512] = ( x[43] );
assign x[513] = ( x[126] );
assign x[514] = ( x[436] );
assign x[515] = ( x[127] );
assign x[516] = ( x[46] );
assign x[517] = ( x[49] );
assign x[518] = ( x[50] );
assign x[519] = ( x[51] );
assign x[520] = ( x[130] );
assign x[521] = ( x[53] );
assign x[522] = ( x[54] );
assign x[523] = ( x[217] );
assign x[524] = ( x[56] );
assign x[525] = ( x[135] );
assign x[526] = ( x[370] );
assign x[527] = ( x[137] );
assign x[528] = ( x[298] );
assign x[529] = ( x[222] );
assign x[530] = ( b & d & e & (~f) & g & h );
assign x[531] = ( x[138] );
assign x[532] = ( x[300] );
assign x[533] = ( x[144] );
assign x[534] = ( x[147] );
assign x[535] = ( x[148] );
assign x[536] = ( x[151] );
assign x[537] = ( x[70] );
assign x[538] = ( x[75] );
assign x[539] = ( x[77] );
assign x[540] = ( b & c & d & (~e) & f );
assign x[541] = ( x[78] );
assign x[542] = ( x[236] );
assign x[543] = ( x[80] );
assign x[544] = ( x[81] );
assign x[545] = ( x[82] );
assign x[546] = ( x[159] );


assign o[1] = |(x[546:468]);



assign x[547] = ( x[389] );
assign x[548] = ( x[471] );
assign x[549] = ( x[390] );
assign x[550] = ( a & (~b) & (~c) & (~d) & (~f) & g & (~h) );
assign x[551] = ( a & b & (~c) & d & (~e) & (~f) & g );
assign x[552] = ( (~a) & b & d & (~e) & f & g & (~h) );
assign x[553] = ( x[2] );
assign x[554] = ( x[86] );
assign x[555] = ( x[320] );
assign x[556] = ( x[87] );
assign x[557] = ( x[165] );
assign x[558] = ( x[89] );
assign x[559] = ( x[90] );
assign x[560] = ( x[250] );
assign x[561] = ( x[482] );
assign x[562] = ( x[175] );
assign x[563] = ( x[257] );
assign x[564] = ( x[99] );
assign x[565] = ( x[489] );
assign x[566] = ( x[100] );
assign x[567] = ( x[263] );
assign x[568] = ( x[27] );
assign x[569] = ( x[266] );
assign x[570] = ( x[28] );
assign x[571] = ( x[187] );
assign x[572] = ( (~a) & c & e & (~f) & g & h );
assign x[573] = ( x[32] );
assign x[574] = ( (~b) & c & (~d) & (~e) & f & g );
assign x[575] = ( (~b) & (~d) & (~e) & (~f) & (~g) & h );
assign x[576] = ( (~a) & c & d & e & f & (~g) );
assign x[577] = ( (~b) & (~c) & d & f & g & (~h) );
assign x[578] = ( a & (~c) & d & f & (~g) & h );
assign x[579] = ( x[196] );
assign x[580] = ( x[111] );
assign x[581] = ( x[112] );
assign x[582] = ( x[281] );
assign x[583] = ( x[36] );
assign x[584] = ( x[282] );
assign x[585] = ( x[357] );
assign x[586] = ( x[283] );
assign x[587] = ( x[37] );
assign x[588] = ( x[287] );
assign x[589] = ( x[118] );
assign x[590] = ( x[41] );
assign x[591] = ( x[44] );
assign x[592] = ( x[436] );
assign x[593] = ( x[210] );
assign x[594] = ( x[46] );
assign x[595] = ( x[50] );
assign x[596] = ( x[51] );
assign x[597] = ( x[130] );
assign x[598] = ( x[131] );
assign x[599] = ( x[53] );
assign x[600] = ( x[54] );
assign x[601] = ( x[217] );
assign x[602] = ( x[55] );
assign x[603] = ( x[56] );
assign x[604] = ( x[371] );
assign x[605] = ( x[220] );
assign x[606] = ( x[530] );
assign x[607] = ( x[58] );
assign x[608] = ( x[372] );
assign x[609] = ( x[59] );
assign x[610] = ( x[140] );
assign x[611] = ( x[141] );
assign x[612] = ( x[142] );
assign x[613] = ( x[65] );
assign x[614] = ( x[144] );
assign x[615] = ( x[147] );
assign x[616] = ( x[69] );
assign x[617] = ( x[74] );
assign x[618] = ( x[236] );
assign x[619] = ( x[80] );
assign x[620] = ( x[82] );


assign o[0] = |(x[620:547]);


endmodule
